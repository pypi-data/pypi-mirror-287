// GENERATE INPLACE BEGIN fileheader() =========================================
//
// Module:     glbl.clk_gate
// Data Model: glbl.clk_gate.ClkGateMod
//
// GENERATE INPLACE END fileheader =============================================

// GENERATE INPLACE BEGIN header() =============================================
`begin_keywords "1800-2009"
`default_nettype none  // implicit wires are forbidden
// GENERATE INPLACE END header =================================================

// GENERATE INPLACE BEGIN beginmod() ===========================================
module clk_gate ( // glbl.clk_gate.ClkGateMod
  input  logic clk_i,
  output logic clk_o,
  input  logic ena_i
);
// GENERATE INPLACE END beginmod ===============================================

    // GENERATE INPLACE BEGIN logic() ==========================================
    // GENERATE INPLACE END logic ==============================================

// GENERATE INPLACE BEGIN endmod() =============================================
endmodule // clk_gate
// GENERATE INPLACE END endmod =================================================

// GENERATE INPLACE BEGIN footer() =============================================
`default_nettype wire
`end_keywords
// GENERATE INPLACE END footer =================================================
