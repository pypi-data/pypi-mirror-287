// GENERATE INPLACE BEGIN fileheader()
// GENERATE INPLACE END fileheader

// GENERATE INPLACE BEGIN header()
// GENERATE INPLACE END header

// GENERATE INPLACE BEGIN beginmod()
// GENERATE INPLACE END beginmod

    // GENERATE INPLACE BEGIN logic()
    // GENERATE INPLACE END logic

// GENERATE INPLACE BEGIN endmod()
// GENERATE INPLACE END endmod

// GENERATE INPLACE BEGIN footer()
// GENERATE INPLACE END footer
